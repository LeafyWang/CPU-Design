//Subject:     CO project 2 - Decoder
//--------------------------------------------------------------------------------
//Version:     1
//--------------------------------------------------------------------------------
//Writer:      
//----------------------------------------------
//Date:        
//----------------------------------------------
//Description: 
//--------------------------------------------------------------------------------

module Decoder(
    instr_op_i,
	RegWrite_o,
	ALU_op_o,
	ALUSrc_o,
	RegDst_o,
	Branch_o
	);
     
//I/O ports
input  [6-1:0] instr_op_i;

output         RegWrite_o;
output [3-1:0] ALU_op_o;
output         ALUSrc_o;
output         RegDst_o;
output         Branch_o;
 
//Internal Signals
reg    [3-1:0] ALU_op_o;
reg            ALUSrc_o;
reg            RegWrite_o;
reg            RegDst_o;
reg            Branch_o;

//Parameter


//Main function
always @(*) begin
case(instr_op_i)
	0: begin ALU_op_o = 3'b010 ; ALUSrc_o = 0;RegWrite_o = 1; RegDst_o = 1;Branch_o = 0; end//add,sub,and,or,slt,sll,srlv
	4: begin ALU_op_o = 3'b001 ; ALUSrc_o = 0;RegWrite_o = 0; RegDst_o = 0;Branch_o = 1; end//beq
        8: begin ALU_op_o = 3'b100 ; ALUSrc_o = 1;RegWrite_o = 1; RegDst_o = 0;Branch_o = 0; end//addi
	10:begin ALU_op_o = 3'b101 ; ALUSrc_o = 1;RegWrite_o = 1; RegDst_o = 0;Branch_o = 0; end//slti
	15:begin ALU_op_o = 3'b011 ; ALUSrc_o = 1;RegWrite_o = 1; RegDst_o = 0;Branch_o = 0; end//lui
	13:begin ALU_op_o = 3'b000 ; ALUSrc_o = 1;RegWrite_o = 1; RegDst_o = 0;Branch_o = 0; end//ori
	5: begin ALU_op_o = 3'b111 ; ALUSrc_o = 0;RegWrite_o = 0; RegDst_o = 0;Branch_o = 1; end//bne
	default:
		begin ALU_op_o = 3'b000 ;ALUSrc_o = 0; RegWrite_o = 0; RegDst_o = 0; Branch_o = 0;end
endcase
end
endmodule





                    
                    